../main.vhdl