../../rotator/src/signed_shifter.vhdl