../main_inst.vhdl