../../uart/src/uart_rx.vhdl