../../uart/src/uart_tx.vhdl