../../ram/implementation/debounce.vhdl