../../rotator/src/cordic.vhdl