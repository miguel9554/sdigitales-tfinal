../../ram/implementation/hex2led.vhdl