../../ram/implementation/disp_mux.vhdl