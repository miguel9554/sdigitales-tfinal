../../uart/src/uart.vhdl