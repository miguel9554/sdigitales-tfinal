../../vga/implementation/xilinx_dual_port_ram_sync.vhdl