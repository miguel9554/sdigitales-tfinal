../../rotator/src/rz.vhdl