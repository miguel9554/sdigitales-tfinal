../../ram/src/sram_controller.vhdl