../../uart/src/fifo.vhdl