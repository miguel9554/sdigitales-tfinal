../../rotator/src/ry.vhdl