../../rotator/src/rx.vhdl