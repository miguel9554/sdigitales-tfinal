../../uart/src/mod_m_counter.vhdl