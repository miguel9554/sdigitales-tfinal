../../vga/src/vga_sync_unit.vhdl