../../rotator/src/addsub.vhdl