../../rotator/src/cordic_stage.vhdl