library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity angle_table is

	port (
		step	:	in unsigned( 3 downto 0);
		angle	:	out unsigned( 21 downto 0)
	);

end entity angle_table;

architecture behavioral of angle_table is

	constant ADDR_WIDTH:	integer	:= 4;
	constant DATA_WIDTH:	integer	:= 22;

	type rom_type is array ( 0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

	constant STEP2ANGLE_ROM: rom_type := (
		"1011010000000000000000",	-- 45°
		"0110101001000010100111",	-- 26.565051177078°
		"0011100000100101000111",	-- 14.0362434679265°
		"0001110010000000000001",	-- 7.1250163489018°
		"0000111001001110001010",	-- 3.57633437499735°
		"0000011100101000110111",	-- 1.78991060824607°
		"0000001110010100101010",	-- 0.895173710211074°
		"0000000111001010010110",	-- 0.447614170860553°
		"0000000011100101001011",	-- 0.223810500368538°
		"0000000001110010100101",	-- 0.111905677066207°
		"0000000000111001010010",	-- 0.055952891893804°
		"0000000000011100101001",	-- 0.027976452617004°
		"0000000000001110010100",	-- 0.013988227142265°
		"0000000000000111001010",	-- 0.006994113675353°
		"0000000000000011100101",	-- 0.003497056850704°
		"0000000000000001110010"	-- 0.00174852842698°
	);

begin

	angle	<=	unsigned(STEP2ANGLE_ROM(to_integer(step)));

end architecture behavioral;