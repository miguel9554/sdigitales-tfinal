../../rotator/src/rotator.vhdl